library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.math_real.all; -- for real numbers

package coefficients is
type coefficients_type is array(0 to 17*4-1) of real;
constant coefficients_250mm_matrix: coefficients_type := (
-- ST matrix 4x4
  0.9966071  ,  1.091514e-2, -2.083274e-3,  3.190145e-4, -- 0*4+
 -0.5563044  ,  0.9438768  , -0.8324718  ,  5.064701e-2, -- 1*4+
  2.153176e-2,  2.126763e-3,  0.7508714  ,  8.221888e-3, -- 2*4+
  3.335013   ,  0.3376467  ,-39.12762    ,  0.4347564  , -- 3*4+
-- PR matrix 1x4
  5.476107e-3,  1.388776   ,  0.2275968  , 35.79262    , -- 4*4+
others => 0.0 -- 5*4+ .. 16*4+ Z0=5*4 and Z1=11*4 variable area
);
-- microcode to calculate one step (ST transposed)
--                            A  = 0  , B = M[0+4*4], C = YP
-- Z0[0]  =   PR[0] * YP      A += B*C, B = M[0+0*4], C = M[0+11*4]
-- Z0[0] += ST[0,0] * Z1[0]   A += B*C, B = M[1+0*4], C = M[1+11*4]
-- Z0[0] += ST[0,1] * Z1[1]   A += B*C, B = M[2+0*4], C = M[2+11*4]
-- Z0[0] += ST[0,2] * Z1[2]   A += B*C, B = M[3+0*4], C = M[3+11*4]
-- Z0[0] += ST[0,3] * Z1[3]   M[0+5*4] = A
--                            A  = 0  , B = M[1+4*4], C = YP
-- Z0[1]  =   PR[1] * YP      A += B*C, B = M[0+1*4], C = M[0+11*4]
-- Z0[1] += ST[1,0] * Z1[0]   A += B*C, B = M[1+1*4], C = M[1+11*4]
-- Z0[1] += ST[1,1] * Z1[1]   A += B*C, B = M[2+1*4], C = M[2+11*4]
-- Z0[1] += ST[1,2] * Z1[2]   A += B*C, B = M[3+1*4], C = M[3+11*4]
-- Z0[1] += ST[1,3] * Z1[3]   M[1+5*4] = A
--                            A  = 0  , B = M[2+4*4], C = YP
-- Z0[2]  =   PR[2] * YP      A += B*C, B = M[0+2*4], C = M[0+11*4]
-- Z0[2] += ST[2,0] * Z1[0]   A += B*C, B = M[1+2*4], C = M[1+11*4]
-- Z0[2] += ST[2,1] * Z1[1]   A += B*C, B = M[2+2*4], C = M[2+11*4]
-- Z0[2] += ST[2,2] * Z1[2]   A += B*C, B = M[3+2*4], C = M[3+11*4]
-- Z0[2] += ST[2,3] * Z1[3]   M[2+5*4] = A
--                            A  = 0  , B = M[3+4*4], C = YP
-- Z0[3]  =   PR[3] * YP      A += B*C, B = M[0+3*4], C = M[0+11*4]
-- Z0[3] += ST[3,0] * Z1[0]   A += B*C, B = M[1+3*4], C = M[1+11*4]
-- Z0[3] += ST[3,1] * Z1[1]   A += B*C, B = M[2+3*4], C = M[2+11*4]
-- Z0[3] += ST[3,2] * Z1[2]   A += B*C, B = M[3+3*4], C = M[3+11*4]
-- Z0[3] += ST[3,3] * Z1[3]   M[3+5*4] = A
--                            A  = 0  , B = M[0+4*4], C = YP
-- Z1[0]  =   PR[0] * YP      A += B*C, B = M[0+0*4], C = M[0+5*4]
-- Z1[0] += ST[0,0] * Z0[0]   A += B*C, B = M[1+0*4], C = M[1+5*4]
-- Z1[0] += ST[0,1] * Z0[1]   A += B*C, B = M[2+0*4], C = M[2+5*4]
-- Z1[0] += ST[0,2] * Z0[2]   A += B*C, B = M[3+0*4], C = M[3+5*4]
-- Z1[0] += ST[0,3] * Z0[3]   M[0+11*4] = A
--                            A  = 0  , B = M[1+4*4], C = YP
-- Z1[1]  =   PR[1] * YP      A += B*C, B = M[0+1*4], C = M[0+5*4]
-- Z1[1] += ST[1,0] * Z0[0]   A += B*C, B = M[1+1*4], C = M[1+5*4]
-- Z1[1] += ST[1,1] * Z0[1]   A += B*C, B = M[2+1*4], C = M[2+5*4]
-- Z1[1] += ST[1,2] * Z0[2]   A += B*C, B = M[3+1*4], C = M[3+5*4]
-- Z1[1] += ST[1,3] * Z0[3]   M[1+11*4] = A
--                            A  = 0  , B = M[2+4*4], C = YP
-- Z1[2]  =   PR[2] * YP      A += B*C, B = M[0+2*4], C = M[0+5*4]
-- Z1[2] += ST[2,0] * Z0[0]   A += B*C, B = M[1+2*4], C = M[1+5*4]
-- Z1[2] += ST[2,1] * Z0[1]   A += B*C, B = M[2+2*4], C = M[2+5*4]
-- Z1[2] += ST[2,2] * Z0[2]   A += B*C, B = M[3+2*4], C = M[3+5*4]
-- Z1[2] += ST[2,3] * Z0[3]   M[2+11*4] = A
--                            A  = 0  , B = M[3+4*4], C = YP
-- Z1[3]  =   PR[3] * YP      A += B*C, B = M[0+3*4], C = M[0+5*4]
-- Z1[3] += ST[3,0] * Z0[0]   A += B*C, B = M[1+3*4], C = M[1+5*4]
-- Z1[3] += ST[3,1] * Z0[1]   A += B*C, B = M[2+3*4], C = M[2+5*4]
-- Z1[3] += ST[3,2] * Z0[2]   A += B*C, B = M[3+3*4], C = M[3+5*4]
-- Z1[3] += ST[3,3] * Z0[3]   M[3+11*4] = A
end coefficients;
