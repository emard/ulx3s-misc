package blinkpkg is
        constant c_blink_bits : natural := 25;
end;
