module top_checkered
(
    input  wire clk_25mhz,
    input  wire [6:0] btn,
    output wire [7:0] led,
    output wire oled_csn,
    output wire oled_clk,
    output wire oled_mosi,
    output wire oled_dc,
    output wire oled_resn,
    output wire wifi_gpio0
);
    assign wifi_gpio0 = btn[0];

    wire clk, locked;
    pll
    pll_inst
    (
        .clki(clk_25mhz),
        .clko(clk), // 12.5 MHz
        .locked(locked)
    );

    wire [6:0] x;
    wire [5:0] y;
    //                 checkered      red     green   blue      red     green   blue
    wire [7:0] color = x[3] ^ y[3] ? {x[6:4], x[6:4], 2'b00} : {y[5:3], 3'b000, 2'b00};

    oled_init
    #(
        .C_init_file("oled_init.mem")
    )
    oled_init_inst
    (
        .clk(clk),
        .x(x),
        .y(y),
        .color(color),
        .oled_csn(oled_csn),
        .oled_clk(oled_clk),
        .oled_mosi(oled_mosi),
        .oled_dc(oled_dc),
        .oled_resn(oled_resn)
    );

endmodule
